configuration tb_meter_cfg of tb_meter is
    for tb
    end for;
  end tb_meter_cfg;
