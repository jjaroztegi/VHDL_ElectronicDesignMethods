configuration tb_div_cfg of tb_div is
    for tb
    end for;
  end tb_div_cfg;