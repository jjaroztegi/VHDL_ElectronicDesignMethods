configuration tb_detector_paridad_cfg of tb_detector_paridad is
    for tb
    end for;
end tb_detector_paridad_cfg;