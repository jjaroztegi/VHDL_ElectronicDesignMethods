configuration tb_decs2p_cfg of tb_decs2p is
    for tb
    end for;
end tb_decs2p_cfg;
