configuration tb_wavegen_cfg of tb_wavegen is
    for tb
    end for;
  end tb_wavegen_cfg;
